netcdf GLASS20006292355 {
dimensions:
	time = 2693 ;
variables:
	int base_time ;
		base_time:long_name = "sounding launch time" ;
		base_time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		base_time:string = "Fri Jun 30 00:49:09 2000" ;
	float time_offset(time) ;
		time_offset:long_name = "seconds since base_time" ;
		time_offset:units = "seconds" ;
		time_offset:missing_value = -999.f ;
		time_offset:_FillValue = -999.f ;
	double time(time) ;
		time:long_name = "time" ;
		time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		time:missing_value = -999.f ;
		time:_FillValue = -999. ;
	float pres(time) ;
		pres:long_name = "pres" ;
		pres:units = "mb" ;
		pres:missing_value = -999.f ;
		pres:_FillValue = -999.f ;
	float tdry(time) ;
		tdry:long_name = "tdry" ;
		tdry:units = "deg C" ;
		tdry:missing_value = -999.f ;
		tdry:_FillValue = -999.f ;
	float dp(time) ;
		dp:long_name = "dp" ;
		dp:units = "deg C" ;
		dp:missing_value = -999.f ;
		dp:_FillValue = -999.f ;
	float rh(time) ;
		rh:long_name = "rh" ;
		rh:units = "percent" ;
		rh:missing_value = -999.f ;
		rh:_FillValue = -999.f ;
	float u_wind(time) ;
		u_wind:long_name = "u_wind" ;
		u_wind:units = "m/s" ;
		u_wind:missing_value = -999.f ;
		u_wind:_FillValue = -999.f ;
	float v_wind(time) ;
		v_wind:long_name = "v_wind" ;
		v_wind:units = "m/s" ;
		v_wind:missing_value = -999.f ;
		v_wind:_FillValue = -999.f ;
	float wspd(time) ;
		wspd:long_name = "wspd" ;
		wspd:units = "m/s" ;
		wspd:missing_value = -999.f ;
		wspd:_FillValue = -999.f ;
	float wdir(time) ;
		wdir:long_name = "wdir" ;
		wdir:units = "degree" ;
		wdir:missing_value = -999.f ;
		wdir:_FillValue = -999.f ;
	float dz(time) ;
		dz:long_name = "dz" ;
		dz:units = "m/s" ;
		dz:missing_value = -999.f ;
		dz:_FillValue = -999.f ;
	float range(time) ;
		range:long_name = "range" ;
		range:units = "km" ;
		range:missing_value = -999.f ;
		range:_FillValue = -999.f ;
	float qp(time) ;
		qp:long_name = "qp" ;
		qp:units = "mb" ;
		qp:missing_value = -999.f ;
		qp:_FillValue = -999.f ;
	float qt(time) ;
		qt:long_name = "qt" ;
		qt:units = "deg C" ;
		qt:missing_value = -999.f ;
		qt:_FillValue = -999.f ;
	float qrh(time) ;
		qrh:long_name = "qrh" ;
		qrh:units = "percent" ;
		qrh:missing_value = -999.f ;
		qrh:_FillValue = -999.f ;
	float qu(time) ;
		qu:long_name = "qu" ;
		qu:units = "m/s" ;
		qu:missing_value = -999.f ;
		qu:_FillValue = -999.f ;
	float qv(time) ;
		qv:long_name = "qv" ;
		qv:units = "m/s" ;
		qv:missing_value = -999.f ;
		qv:_FillValue = -999.f ;
	float qwind(time) ;
		qwind:long_name = "qwind" ;
		qwind:units = "m/s" ;
		qwind:missing_value = -999.f ;
		qwind:_FillValue = -999.f ;
	float mr(time) ;
		mr:long_name = "mr" ;
		mr:units = "g/kg" ;
		mr:missing_value = -999.f ;
		mr:_FillValue = -999.f ;
	float vt(time) ;
		vt:long_name = "vt" ;
		vt:units = "deg C" ;
		vt:missing_value = -999.f ;
		vt:_FillValue = -999.f ;
	float theta(time) ;
		theta:long_name = "theta" ;
		theta:units = "deg K" ;
		theta:missing_value = -999.f ;
		theta:_FillValue = -999.f ;
	float theta_e(time) ;
		theta_e:long_name = "theta_e" ;
		theta_e:units = "deg K" ;
		theta_e:missing_value = -999.f ;
		theta_e:_FillValue = -999.f ;
	float theta_v(time) ;
		theta_v:long_name = "theta_v" ;
		theta_v:units = "deg K" ;
		theta_v:missing_value = -999.f ;
		theta_v:_FillValue = -999.f ;
	float lat(time) ;
		lat:long_name = "north latitude" ;
		lat:units = "degrees" ;
		lat:missing_value = -999.f ;
		lat:_FillValue = -999.f ;
		lat:valid_range = -90.f, 90.f ;
	float lon(time) ;
		lon:long_name = "east longitude" ;
		lon:units = "degrees" ;
		lon:missing_value = -999.f ;
		lon:_FillValue = -999.f ;
		lon:valid_range = -180.f, 180.f ;
	float alt(time) ;
		alt:long_name = "altitude" ;
		alt:units = "meters" ;
		alt:missing_value = -999.f ;
		alt:_FillValue = -999.f ;

// global attributes:
		:bad_value_flag = -999.f ;
		:zebra_platform = "class" ;
		:history = "ClassNcFile" ;
		:AvapsEditorVersion = "2.2.2" ;
		:SoundingDescription = "D200006292355.st1 Version:       STEPS Mobile 1, GLASS 2.01\r  " ;
		:ACagency = "AF001" ;
		:ACtype = "0" ;
		:AbrHdrOvr = "0" ;
		:BaudRateIndex = "2" ;
		:CommPortIndex = "0" ;
		:IcaoIndex = "1" ;
		:MissionId = "TRAIN" ;
		:MissionStorm = "WXWXA" ;
		:OptIcao = "W" ;
		:OptionAutoFile = "1" ;
		:OptionBSN = "99999" ;
		:OptionCallSign = "CALL" ;
		:OptionChuteArea = "676" ;
		:OptionDoLevels = "1" ;
		:OptionDoQC = "1" ;
		:OptionDoWMO = "1" ;
		:OptionDropSondeMass = "395" ;
		:OptionPosInterpSpan = "60" ;
		:OptionTempMsgType = "2" ;
		:PresBuddySlope = "2" ;
		:PresOffset = "0" ;
		:PresOutlier = "10" ;
		:PresQCDev = "3" ;
		:PresQCWL = "60" ;
		:PresSmoothWL = "60" ;
		:QCSaveDir = "H:\\steps" ;
		:RHBuddySlope = "20" ;
		:RHOffset = "0" ;
		:RHOutlier = "10" ;
		:RHQCDev = "3" ;
		:RHQCWL = "60" ;
		:RHSmoothWL = "60" ;
		:RawSaveDir = "6" ;
		:SfcAltUnknown = "0" ;
		:SfcAltitude = "955.1" ;
		:TdryBuddySlope = "3" ;
		:TdryDynCor = "1" ;
		:TdryOffset = "0" ;
		:TdryOutlier = "10" ;
		:TdryQCDev = "3" ;
		:TdryQCWL = "60" ;
		:TdrySmoothWL = "60" ;
		:WindBuddySlope = "5" ;
		:WindDynCor = "1" ;
		:WindOutlier = "10" ;
		:WindQCDev = "3" ;
		:WindQCWL = "10" ;
		:WindSats = "3" ;
		:WindSmoothWL = "10" ;
		:WindVVdelta = "2.5" ;
		:WmoSaveDir = "C:\\" ;
		:excludeAbrHdr = "0" ;
data:

 time = 962347748, 962347749, 962347750, 962347751, 962347752, 962347753, 
    962347754, 962347755, 962347756, 962347757, 962347758, 962347759, 
    962347760, 962347761, 962347762, 962347763, 962347764, 962347765, 
    962347766, 962347767, 962347768, 962347769, 962347770, 962347771, 
    962347772, 962347773, 962347774, 962347775, 962347776, 962347777, 
    962347778, 962347779, 962347780, 962347781, 962347782, 962347783, 
    962347784, 962347785, 962347786, 962347787, 962347788, 962347789, 
    962347790, 962347791, 962347792, 962347793, 962347794, 962347795, 
    962347796, 962347797, 962347798, 962347799, 962347800, 962347801, 
    962347802, 962347803, 962347804, 962347805, 962347806, 962347807, 
    962347808.1, 962347809.1, 962347810.1, 962347811.1, 962347812.1, 
    962347813.1, 962347814.1, 962347815.1, 962347816.1, 962347817.1, 
    962347818.1, 962347819.1, 962347820.1, 962347821.1, 962347822.1, 
    962347823.1, 962347824.1, 962347825.1, 962347826.1, 962347827.1, 
    962347828.1, 962347829.1, 962347830.1, 962347831.1, 962347832.1, 
    962347833.1, 962347834.1, 962347835.1, 962347836.1, 962347837.1, 
    962347838.1, 962347839.1, 962347840.1, 962347841.1, 962347842.1, 
    962347843.1, 962347844.1, 962347845.1, 962347846.1, 962347847.1, 
    962347848.1, 962347849.1, 962347850.1, 962347851.1, 962347852.1, 
    962347853.1, 962347854.1, 962347855.1, 962347856.1, 962347857.1, 
    962347858.1, 962347859.1, 962347860.1, 962347861.1, 962347862.1, 
    962347863.1, 962347864.1, 962347865.1, 962347866.1, 962347867.1, 
    962347868.1, 962347869.1, 962347870.1, 962347871.1, 962347872.1, 
    962347873.1, 962347874.1, 962347875.1, 962347876.1, 962347877.1, 
    962347878.1, 962347879.1, 962347880.1, 962347881.1, 962347882.1, 
    962347883.1, 962347884.1, 962347885.1, 962347886.1, 962347887.1, 
    962347888.1, 962347889.1, 962347890.1, 962347891.1, 962347892.1, 
    962347893.1, 962347894.1, 962347895.1, 962347896.1, 962347897.1, 
    962347898.1, 962347899.1, 962347900.1, 962347901.1, 962347902.1, 
    962347903.1, 962347904.1, 962347905.1, 962347906.1, 962347907.2, 
    962347908.2, 962347909.2, 962347910.2, 962347911.2, 962347912.2, 
    962347913.2, 962347914.2, 962347915.2, 962347916.2, 962347917.2, 
    962347918.2, 962347919.2, 962347920.2, 962347921.2, 962347922.2, 
    962347923.2, 962347924.2, 962347925.2, 962347926.2, 962347927.2, 
    962347928.2, 962347929.2, 962347930.2, 962347931.2, 962347932.2, 
    962347933.2, 962347934.2, 962347935.2, 962347936.2, 962347937.2, 
    962347938.2, 962347939.2, 962347940.2, 962347941.2, 962347942.2, 
    962347943.2, 962347944.2, 962347945.2, 962347946.2, 962347947.2, 
    962347948.2, 962347949.2, 962347950.2, 962347951.2, 962347952.2, 
    962347953.2, 962347954.2, 962347955.2, 962347956.2, 962347957.2, 
    962347958.2, 962347959.2, 962347960.2, 962347961.2, 962347962.2, 
    962347963.2, 962347964.2, 962347965.2, 962347966.2, 962347967.2, 
    962347968.2, 962347969.2, 962347970.2, 962347971.2, 962347972.2, 
    962347973.2, 962347974.2, 962347975.2, 962347976.2, 962347977.2, 
    962347978.2, 962347979.2, 962347980.2, 962347981.2, 962347982.2, 
    962347983.2, 962347984.2, 962347985.2, 962347986.2, 962347987.2, 
    962347988.2, 962347989.2, 962347990.2, 962347991.2, 962347992.2, 
    962347993.2, 962347994.2, 962347995.2, 962347996.2, 962347997.2, 
    962347998.2, 962347999.2, 962348000.2, 962348001.2, 962348002.2, 
    962348003.2, 962348004.2, 962348005.2, 962348006.2, 962348007.2, 
    962348008.2, 962348009.2, 962348010.2, 962348011.3, 962348012.3, 
    962348013.3, 962348014.3, 962348015.3, 962348016.3, 962348017.3, 
    962348018.3, 962348019.3, 962348020.3, 962348021.3, 962348022.3, 
    962348023.3, 962348024.3, 962348025.3, 962348026.3, 962348027.3, 
    962348028.3, 962348029.3, 962348030.3, 962348031.3, 962348032.3, 
    962348033.3, 962348034.3, 962348035.3, 962348036.3, 962348037.3, 
    962348038.3, 962348039.3, 962348040.3, 962348041.3, 962348042.3, 
    962348043.3, 962348044.3, 962348045.3, 962348046.3, 962348047.3, 
    962348048.3, 962348049.3, 962348050.3, 962348051.3, 962348052.3, 
    962348053.3, 962348054.3, 962348055.3, 962348056.3, 962348057.3, 
    962348058.3, 962348059.3, 962348060.3, 962348061.3, 962348062.3, 
    962348063.3, 962348064.3, 962348065.3, 962348066.3, 962348067.3, 
    962348068.3, 962348069.3, 962348070.3, 962348071.3, 962348072.3, 
    962348073.3, 962348074.3, 962348075.3, 962348076.3, 962348077.3, 
    962348078.3, 962348079.3, 962348080.3, 962348081.3, 962348082.3, 
    962348083.3, 962348084.3, 962348085.3, 962348086.3, 962348087.3, 
    962348088.3, 962348089.3, 962348090.3, 962348091.3, 962348092.3, 
    962348093.3, 962348094.3, 962348095.3, 962348096.3, 962348097.3, 
    962348098.3, 962348099.3, 962348100.3, 962348101.3, 962348102.3, 
    962348103.3, 962348104.3, 962348105.3, 962348106.3, 962348107.3, 
    962348108.3, 962348109.3, 962348110.3, 962348111.3, 962348112.3, 
    962348113.4, 962348114.4, 962348115.4, 962348116.4, 962348117.4, 
    962348118.4, 962348119.4, 962348120.4, 962348121.4, 962348122.4, 
    962348123.4, 962348124.4, 962348125.4, 962348126.4, 962348127.4, 
    962348128.4, 962348129.4, 962348130.4, 962348131.4, 962348132.4, 
    962348133.4, 962348134.4, 962348135.4, 962348136.4, 962348137.4, 
    962348138.4, 962348139.4, 962348140.4, 962348141.4, 962348142.4, 
    962348143.4, 962348144.4, 962348145.4, 962348146.4, 962348147.4, 
    962348148.4, 962348149.4, 962348150.4, 962348151.4, 962348152.4, 
    962348153.4, 962348154.4, 962348155.4, 962348156.4, 962348157.4, 
    962348158.4, 962348159.4, 962348160.4, 962348161.4, 962348162.4, 
    962348163.4, 962348164.4, 962348165.4, 962348166.4, 962348167.4, 
    962348168.4, 962348169.4, 962348170.4, 962348171.4, 962348172.4, 
    962348173.4, 962348174.4, 962348175.4, 962348176.4, 962348177.4, 
    962348178.4, 962348179.4, 962348180.4, 962348181.4, 962348182.4, 
    962348183.4, 962348184.4, 962348185.4, 962348186.4, 962348187.4, 
    962348188.4, 962348189.4, 962348190.4, 962348191.4, 962348192.4, 
    962348193.4, 962348194.4, 962348195.4, 962348196.4, 962348197.4, 
    962348198.4, 962348199.4, 962348200.4, 962348201.4, 962348202.4, 
    962348203.4, 962348204.4, 962348205.5, 962348206.5, 962348207.5, 
    962348208.5, 962348209.5, 962348210.5, 962348211.5, 962348212.5, 
    962348213.5, 962348214.5, 962348215.5, 962348216.5, 962348217.5, 
    962348218.5, 962348219.5, 962348220.5, 962348221.5, 962348222.5, 
    962348223.5, 962348224.5, 962348225.5, 962348226.5, 962348227.5, 
    962348228.5, 962348229.5, 962348230.5, 962348231.5, 962348232.5, 
    962348233.5, 962348234.5, 962348235.5, 962348236.5, 962348237.5, 
    962348238.5, 962348239.5, 962348240.5, 962348241.5, 962348242.5, 
    962348243.5, 962348244.5, 962348245.5, 962348246.5, 962348247.5, 
    962348248.5, 962348249.5, 962348250.5, 962348251.5, 962348252.5, 
    962348253.5, 962348254.5, 962348255.5, 962348256.5, 962348257.5, 
    962348258.5, 962348259.5, 962348260.5, 962348261.5, 962348262.5, 
    962348263.5, 962348264.5, 962348265.5, 962348266.5, 962348267.5, 
    962348268.5, 962348269.5, 962348270.5, 962348271.5, 962348272.5, 
    962348273.5, 962348274.5, 962348275.5, 962348276.5, 962348277.5, 
    962348278.5, 962348279.5, 962348280.5, 962348281.5, 962348282.5, 
    962348283.5, 962348284.5, 962348285.5, 962348286.5, 962348287.5, 
    962348288.5, 962348289.5, 962348290.5, 962348291.5, 962348292.5, 
    962348293.5, 962348294.5, 962348295.5, 962348296.5, 962348297.5, 
    962348298.5, 962348299.5, 962348300.5, 962348301.5, 962348302.5, 
    962348303.5, 962348304.5, 962348305.5, 962348306.5, 962348307.5, 
    962348308.5, 962348309.5, 962348310.5, 962348311.5, 962348312.5, 
    962348313.5, 962348314.5, 962348315.5, 962348316.5, 962348317.6, 
    962348318.6, 962348319.6, 962348320.6, 962348321.6, 962348322.6, 
    962348323.6, 962348324.6, 962348325.6, 962348326.6, 962348327.6, 
    962348328.6, 962348329.6, 962348330.6, 962348331.6, 962348332.6, 
    962348333.6, 962348334.6, 962348335.6, 962348336.6, 962348337.6, 
    962348338.6, 962348339.6, 962348340.6, 962348341.6, 962348342.6, 
    962348343.6, 962348344.6, 962348345.6, 962348346.6, 962348347.6, 
    962348348.6, 962348349.6, 962348350.6, 962348351.6, 962348352.6, 
    962348353.6, 962348354.6, 962348355.6, 962348356.6, 962348357.6, 
    962348358.6, 962348359.6, 962348360.6, 962348361.6, 962348362.6, 
    962348363.6, 962348364.6, 962348365.6, 962348366.6, 962348367.6, 
    962348368.6, 962348369.6, 962348370.6, 962348371.6, 962348372.6, 
    962348373.6, 962348374.6, 962348375.6, 962348376.6, 962348377.6, 
    962348378.6, 962348379.6, 962348380.6, 962348381.6, 962348382.6, 
    962348383.6, 962348384.6, 962348385.6, 962348386.6, 962348387.6, 
    962348388.6, 962348389.6, 962348390.6, 962348391.6, 962348392.6, 
    962348393.6, 962348394.6, 962348395.6, 962348396.6, 962348397.6, 
    962348398.6, 962348399.6, 962348400.6, 962348401.6, 962348402.6, 
    962348403.6, 962348404.6, 962348405.6, 962348406.6, 962348407.6, 
    962348408.6, 962348409.7, 962348410.7, 962348411.7, 962348412.7, 
    962348413.7, 962348414.7, 962348415.7, 962348416.7, 962348417.7, 
    962348418.7, 962348419.7, 962348420.7, 962348421.7, 962348422.7, 
    962348423.7, 962348424.7, 962348425.7, 962348426.7, 962348427.7, 
    962348428.7, 962348429.7, 962348430.7, 962348431.7, 962348432.7, 
    962348433.7, 962348434.7, 962348435.7, 962348436.7, 962348437.7, 
    962348438.7, 962348439.7, 962348440.7, 962348441.7, 962348442.7, 
    962348443.7, 962348444.7, 962348445.7, 962348446.7, 962348447.7, 
    962348448.7, 962348449.7, 962348450.7, 962348451.7, 962348452.7, 
    962348453.7, 962348454.7, 962348455.7, 962348456.7, 962348457.7, 
    962348458.7, 962348459.7, 962348460.7, 962348461.7, 962348462.7, 
    962348463.7, 962348464.7, 962348465.7, 962348466.7, 962348467.7, 
    962348468.7, 962348469.7, 962348470.7, 962348471.7, 962348472.7, 
    962348473.7, 962348474.7, 962348475.7, 962348476.7, 962348477.7, 
    962348478.7, 962348479.7, 962348480.7, 962348481.7, 962348482.7, 
    962348483.7, 962348484.7, 962348485.7, 962348486.7, 962348487.7, 
    962348488.7, 962348489.7, 962348490.7, 962348491.7, 962348492.7, 
    962348493.7, 962348494.7, 962348495.7, 962348496.7, 962348497.7, 
    962348498.7, 962348499.7, 962348500.7, 962348501.7, 962348502.7, 
    962348503.7, 962348504.7, 962348505.7, 962348506.7, 962348507.7, 
    962348508.7, 962348509.7, 962348510.7, 962348511.8, 962348512.8, 
    962348513.8, 962348514.8, 962348515.8, 962348516.8, 962348517.8, 
    962348518.8, 962348519.8, 962348520.8, 962348521.8, 962348522.8, 
    962348523.8, 962348524.8, 962348525.8, 962348526.8, 962348527.8, 
    962348528.8, 962348529.8, 962348530.8, 962348531.8, 962348532.8, 
    962348533.8, 962348534.8, 962348535.8, 962348536.8, 962348537.8, 
    962348538.8, 962348539.8, 962348540.8, 962348541.8, 962348542.8, 
    962348543.8, 962348544.8, 962348545.8, 962348546.8, 962348547.8, 
    962348548.8, 962348549.8, 962348550.8, 962348551.8, 962348552.8, 
    962348553.8, 962348554.8, 962348555.8, 962348556.8, 962348557.8, 
    962348558.8, 962348559.8, 962348560.8, 962348561.8, 962348562.8, 
    962348563.3, 962348564.3, 962348565.3, 962348566.3, 962348567.3, 
    962348568.3, 962348569.3, 962348570.3, 962348571.3, 962348572.3, 
    962348573.3, 962348574.3, 962348575.3, 962348576.3, 962348577.3, 
    962348578.3, 962348579.3, 962348580.3, 962348581.3, 962348582.3, 
    962348583.3, 962348584.3, 962348585.3, 962348586.3, 962348587.3, 
    962348588.3, 962348589.3, 962348590.3, 962348591.3, 962348592.3, 
    962348593.3, 962348594.3, 962348595.3, 962348596.3, 962348597.3, 
    962348598.3, 962348599.3, 962348600.3, 962348601.3, 962348602.3, 
    962348603.3, 962348604.3, 962348605.3, 962348606.3, 962348607.3, 
    962348608.3, 962348609.3, 962348610.3, 962348611.3, 962348612.3, 
    962348613.4, 962348614.4, 962348615.4, 962348616.4, 962348617.4, 
    962348618.4, 962348619.4, 962348620.4, 962348621.4, 962348622.4, 
    962348623.4, 962348624.4, 962348625.4, 962348626.4, 962348627.4, 
    962348628.4, 962348629.4, 962348630.4, 962348631.4, 962348632.4, 
    962348633.4, 962348634.4, 962348635.4, 962348636.4, 962348637.4, 
    962348638.4, 962348639.4, 962348640.4, 962348641.4, 962348642.4, 
    962348643.4, 962348644.4, 962348645.4, 962348646.4, 962348647.4, 
    962348648.4, 962348649.4, 962348650.4, 962348651.4, 962348652.4, 
    962348653.4, 962348654.4, 962348655.4, 962348656.4, 962348657.4, 
    962348658.4, 962348659.4, 962348660.4, 962348661.4, 962348662.4, 
    962348663.4, 962348664.4, 962348665.4, 962348666.4, 962348667.4, 
    962348668.4, 962348669.4, 962348670.4, 962348671.4, 962348672.4, 
    962348673.4, 962348674.4, 962348675.4, 962348676.4, 962348677.4, 
    962348678.4, 962348679.4, 962348680.4, 962348681.4, 962348682.4, 
    962348683.4, 962348684.4, 962348685.4, 962348686.4, 962348687.4, 
    962348688.4, 962348689.4, 962348690.4, 962348691.4, 962348692.4, 
    962348693.4, 962348694.4, 962348695.4, 962348696.4, 962348697.4, 
    962348698.4, 962348699.4, 962348700.4, 962348701.4, 962348702.4, 
    962348703.4, 962348704.4, 962348705.4, 962348706.4, 962348707.4, 
    962348708.4, 962348709.4, 962348710.4, 962348711.4, 962348712.4, 
    962348713.4, 962348714.4, 962348715.5, 962348716.5, 962348717.5, 
    962348718.5, 962348719.5, 962348720.5, 962348721.5, 962348722.5, 
    962348723.5, 962348724.5, 962348725.5, 962348726.5, 962348727.5, 
    962348728.5, 962348729.5, 962348730.5, 962348731.5, 962348732.5, 
    962348733.5, 962348734.5, 962348735.5, 962348736.5, 962348737.5, 
    962348738.5, 962348739.5, 962348740.5, 962348741.5, 962348742.5, 
    962348743.5, 962348744.5, 962348745.5, 962348746.5, 962348747.5, 
    962348748.5, 962348749.5, 962348750.5, 962348751.5, 962348752.5, 
    962348753.5, 962348754.5, 962348755.5, 962348756, 962348757, 962348758, 
    962348759, 962348760, 962348761, 962348762, 962348763, 962348764, 
    962348765, 962348766, 962348767, 962348768, 962348769, 962348770, 
    962348771, 962348772, 962348773, 962348774, 962348775, 962348776, 
    962348777, 962348778, 962348779, 962348780, 962348781, 962348782, 
    962348783, 962348784, 962348785, 962348786, 962348787, 962348788, 
    962348789, 962348790, 962348791, 962348792, 962348793, 962348794, 
    962348795, 962348796, 962348797, 962348798, 962348799, 962348800, 
    962348801, 962348802, 962348803, 962348804, 962348805, 962348806, 
    962348807, 962348808, 962348809, 962348810, 962348811, 962348812, 
    962348813, 962348814, 962348815, 962348816, 962348817, 962348818, 
    962348819, 962348820, 962348821, 962348822, 962348823, 962348824, 
    962348825, 962348826, 962348827, 962348828.1, 962348829.1, 962348830.1, 
    962348831.1, 962348832.1, 962348833.1, 962348834.1, 962348835.1, 
    962348836.1, 962348837.1, 962348838.1, 962348839.1, 962348840.1, 
    962348841.1, 962348842.1, 962348843.1, 962348844.1, 962348845.1, 
    962348846.1, 962348847.1, 962348848.1, 962348848.6, 962348849.6, 
    962348850.6, 962348851.6, 962348852.6, 962348853.6, 962348854.6, 
    962348855.6, 962348856.6, 962348857.6, 962348858.6, 962348859.6, 
    962348860.6, 962348861.6, 962348862.6, 962348863.6, 962348864.6, 
    962348865.6, 962348866.6, 962348867.6, 962348868.6, 962348869.6, 
    962348870.6, 962348871.6, 962348872.6, 962348873.6, 962348874.6, 
    962348875.6, 962348876.6, 962348877.6, 962348878.6, 962348879.6, 
    962348880.6, 962348881.6, 962348882.6, 962348883.6, 962348884.6, 
    962348885.6, 962348886.6, 962348887.6, 962348888.6, 962348889.6, 
    962348890.6, 962348891.6, 962348892.6, 962348893.6, 962348894.6, 
    962348895.6, 962348896.6, 962348897.6, 962348898.6, 962348899.6, 
    962348900.6, 962348901.6, 962348902.6, 962348903.6, 962348904.6, 
    962348905.6, 962348906.6, 962348907.6, 962348908.6, 962348909.6, 
    962348910.6, 962348911.6, 962348912.6, 962348913.6, 962348914.6, 
    962348915.6, 962348916.6, 962348917.6, 962348918.6, 962348919.6, 
    962348920.6, 962348921.6, 962348922.6, 962348923.6, 962348924.6, 
    962348925.6, 962348926.6, 962348927.6, 962348928.6, 962348929.6, 
    962348930.2, 962348931.2, 962348932.2, 962348933.2, 962348934.2, 
    962348935.2, 962348936.2, 962348937.2, 962348938.2, 962348939.2, 
    962348940.2, 962348941.2, 962348942.2, 962348943.2, 962348944.2, 
    962348945.2, 962348946.2, 962348947.2, 962348948.2, 962348949.2, 
    962348950.2, 962348951.2, 962348952.2, 962348953.2, 962348954.2, 
    962348955.2, 962348956.2, 962348957.2, 962348958.2, 962348959.2, 
    962348960.2, 962348961.2, 962348962.2, 962348963.2, 962348964.2, 
    962348965.2, 962348966.2, 962348967.2, 962348968.2, 962348969.2, 
    962348970.2, 962348971.2, 962348972.2, 962348973.2, 962348974.2, 
    962348975.2, 962348976.2, 962348977.2, 962348978.2, 962348979.2, 
    962348980.2, 962348981.2, 962348982.2, 962348983.2, 962348984.2, 
    962348985.2, 962348986.2, 962348987.2, 962348988.2, 962348989.2, 
    962348990.2, 962348991.2, 962348992.2, 962348993.2, 962348994.2, 
    962348995.2, 962348996.2, 962348997.2, 962348998.2, 962348999.2, 
    962349000.2, 962349001.2, 962349002.2, 962349003.2, 962349004.2, 
    962349005.2, 962349006.2, 962349007.2, 962349008.2, 962349009.2, 
    962349010.2, 962349011.2, 962349011.7, 962349012.7, 962349013.7, 
    962349014.7, 962349015.7, 962349016.7, 962349017.7, 962349018.7, 
    962349019.7, 962349020.7, 962349021.8, 962349022.8, 962349023.8, 
    962349024.8, 962349025.8, 962349026.8, 962349027.8, 962349028.8, 
    962349029.8, 962349030.8, 962349031.8, 962349032.8, 962349033.8, 
    962349034.8, 962349035.8, 962349036.8, 962349037.8, 962349038.8, 
    962349039.8, 962349040.8, 962349041.8, 962349042.8, 962349043.8, 
    962349044.8, 962349045.8, 962349046.8, 962349047.8, 962349048.8, 
    962349049.8, 962349050.8, 962349051.8, 962349052.8, 962349053.8, 
    962349054.8, 962349055.8, 962349056.8, 962349057.8, 962349058.8, 
    962349059.8, 962349060.8, 962349061.8, 962349062.8, 962349063.8, 
    962349064.8, 962349065.8, 962349066.8, 962349067.8, 962349068.8, 
    962349069.8, 962349070.8, 962349071.8, 962349072.3, 962349073.3, 
    962349074.3, 962349075.3, 962349076.3, 962349077.3, 962349078.3, 
    962349079.3, 962349080.3, 962349081.3, 962349082.3, 962349083.3, 
    962349084.3, 962349085.3, 962349086.3, 962349087.3, 962349088.3, 
    962349089.3, 962349090.3, 962349091.3, 962349092.3, 962349093.3, 
    962349094.3, 962349095.3, 962349096.3, 962349097.3, 962349098.3, 
    962349099.3, 962349100.3, 962349101.3, 962349102.3, 962349103.3, 
    962349104.3, 962349105.3, 962349106.3, 962349107.3, 962349108.3, 
    962349109.3, 962349110.3, 962349111.3, 962349112.3, 962349113.3, 
    962349113.8, 962349114.8, 962349115.8, 962349116.8, 962349117.8, 
    962349118.8, 962349119.8, 962349120.8, 962349121.8, 962349122.8, 
    962349123.9, 962349124.9, 962349125.9, 962349126.9, 962349127.9, 
    962349128.9, 962349129.9, 962349130.9, 962349131.9, 962349132.9, 
    962349133.9, 962349134.9, 962349135.9, 962349136.9, 962349137.9, 
    962349138.9, 962349139.9, 962349140.9, 962349141.9, 962349142.9, 
    962349143.9, 962349144.9, 962349145.9, 962349146.9, 962349147.9, 
    962349148.9, 962349149.9, 962349150.9, 962349151.9, 962349152.9, 
    962349153.9, 962349154.9, 962349155.9, 962349156.9, 962349157.9, 
    962349158.9, 962349159.9, 962349160.9, 962349161.9, 962349162.9, 
    962349163.9, 962349164.9, 962349165.9, 962349166.9, 962349167.9, 
    962349168.9, 962349169.9, 962349170.9, 962349171.9, 962349172.9, 
    962349173.9, 962349174.9, 962349175.9, 962349176.9, 962349177.9, 
    962349178.9, 962349179.9, 962349180.9, 962349181.9, 962349182.9, 
    962349183.9, 962349184.9, 962349185.9, 962349186.9, 962349187.9, 
    962349188.9, 962349189.9, 962349190.9, 962349191.9, 962349192.9, 
    962349193.9, 962349194.9, 962349195.9, 962349196.9, 962349197.9, 
    962349198.9, 962349199.9, 962349200.9, 962349201.9, 962349202.9, 
    962349203.9, 962349204.9, 962349205.9, 962349206.9, 962349207.9, 
    962349208.9, 962349209.9, 962349210.9, 962349211.9, 962349212.9, 
    962349213.9, 962349214.9, 962349215.4, 962349216.4, 962349217.4, 
    962349218.4, 962349219.4, 962349220.4, 962349221.4, 962349222.4, 
    962349223.4, 962349224.4, 962349225.5, 962349226.5, 962349227.5, 
    962349228.5, 962349229.5, 962349230.5, 962349231.5, 962349232.5, 
    962349233.5, 962349234.5, 962349235.5, 962349236.5, 962349237.5, 
    962349238.5, 962349239.5, 962349240.5, 962349241.5, 962349242.5, 
    962349243.5, 962349244.5, 962349245.5, 962349246.5, 962349247.5, 
    962349248.5, 962349249.5, 962349250.5, 962349251.5, 962349252.5, 
    962349253.5, 962349254.5, 962349255.5, 962349256.5, 962349257.5, 
    962349258.5, 962349259.5, 962349260.5, 962349261.5, 962349262.5, 
    962349263.5, 962349264.5, 962349265.5, 962349266.5, 962349267.5, 
    962349268.5, 962349269.5, 962349270.5, 962349271.5, 962349272.5, 
    962349273.5, 962349274.5, 962349275.5, 962349276.5, 962349277.5, 
    962349278.5, 962349279.5, 962349280.5, 962349281.5, 962349282.5, 
    962349283.5, 962349284.5, 962349285.5, 962349286.5, 962349287.5, 
    962349288.5, 962349289.5, 962349290.5, 962349291.5, 962349292.5, 
    962349293.5, 962349294.5, 962349295.5, 962349296.5, 962349297, 962349298, 
    962349299, 962349300, 962349301, 962349302, 962349303, 962349304, 
    962349305, 962349306, 962349307, 962349308, 962349309, 962349310, 
    962349311, 962349312, 962349313, 962349314, 962349315, 962349316, 
    962349317, 962349318, 962349319, 962349320, 962349321, 962349322, 
    962349323, 962349324, 962349325, 962349326, 962349327, 962349328, 
    962349329, 962349330, 962349331, 962349332, 962349333, 962349334, 
    962349335, 962349336, 962349337, 962349338.1, 962349339.1, 962349340.1, 
    962349341.1, 962349342.1, 962349343.1, 962349344.1, 962349345.1, 
    962349346.1, 962349347.1, 962349348.1, 962349349.1, 962349350.1, 
    962349351.1, 962349352.1, 962349353.1, 962349354.1, 962349355.1, 
    962349356.1, 962349357.1, 962349358.1, 962349359.1, 962349360.1, 
    962349361.1, 962349362.1, 962349363.1, 962349364.1, 962349365.1, 
    962349366.1, 962349367.1, 962349368.1, 962349369.1, 962349370.1, 
    962349371.1, 962349372.1, 962349373.1, 962349374.1, 962349375.1, 
    962349376.1, 962349377.1, 962349378.1, 962349379.1, 962349380.1, 
    962349381.1, 962349382.1, 962349383.1, 962349384.1, 962349385.1, 
    962349386.1, 962349387.1, 962349388.1, 962349389.1, 962349390.1, 
    962349391.1, 962349392.1, 962349393.1, 962349394.1, 962349395.1, 
    962349396.1, 962349397.1, 962349398.1, 962349399.1, 962349400.1, 
    962349401.1, 962349402.1, 962349403.1, 962349404.1, 962349405.1, 
    962349406.1, 962349407.1, 962349408.1, 962349409.1, 962349410.1, 
    962349411.1, 962349412.1, 962349413.1, 962349414.1, 962349415.1, 
    962349416.1, 962349417.1, 962349418.1, 962349419.1, 962349420.1, 
    962349421.1, 962349422.1, 962349423.1, 962349424.1, 962349425.1, 
    962349426.1, 962349427.1, 962349428.1, 962349429.1, 962349430.1, 
    962349431.1, 962349432.1, 962349433.1, 962349434.1, 962349435.1, 
    962349436.1, 962349437.1, 962349438.1, 962349439.1, 962349440.2, 
    962349441.2, 962349442.2, 962349443.2, 962349444.2, 962349445.2, 
    962349446.2, 962349447.2, 962349448.2, 962349449.2, 962349450.2, 
    962349451.2, 962349452.2, 962349453.2, 962349454.2, 962349455.2, 
    962349456.2, 962349457.2, 962349458.2, 962349459.2, 962349460.2, 
    962349461.2, 962349462.2, 962349463.2, 962349464.2, 962349465.2, 
    962349466.2, 962349467.2, 962349468.2, 962349469.2, 962349470.2, 
    962349471.2, 962349472.2, 962349473.2, 962349474.2, 962349475.2, 
    962349476.2, 962349477.2, 962349478.2, 962349479.2, 962349480.2, 
    962349481.2, 962349482.2, 962349483.2, 962349484.2, 962349485.2, 
    962349486.2, 962349487.2, 962349488.2, 962349489.2, 962349490.2, 
    962349491.2, 962349492.2, 962349493.2, 962349494.2, 962349495.2, 
    962349496.2, 962349497.2, 962349498.2, 962349499.2, 962349500.2, 
    962349501.2, 962349502.2, 962349503.2, 962349504.2, 962349505.2, 
    962349506.2, 962349507.2, 962349508.2, 962349509.2, 962349510.2, 
    962349511.2, 962349512.2, 962349512.7, 962349513.7, 962349514.7, 
    962349515.7, 962349516.7, 962349517.7, 962349518.7, 962349519.7, 
    962349520.7, 962349521.7, 962349522.2, 962349523.2, 962349524.2, 
    962349525.2, 962349526.2, 962349527.2, 962349528.2, 962349529.2, 
    962349530.2, 962349531.2, 962349532.3, 962349533.3, 962349534.3, 
    962349535.3, 962349536.3, 962349537.3, 962349538.3, 962349539.3, 
    962349540.3, 962349541.3, 962349542.3, 962349543.3, 962349544.3, 
    962349545.3, 962349546.3, 962349547.3, 962349548.3, 962349549.3, 
    962349550.3, 962349551.3, 962349551.8, 962349552.8, 962349553.8, 
    962349554.8, 962349555.8, 962349556.8, 962349557.8, 962349558.8, 
    962349559.8, 962349560.8, 962349561.8, 962349562.3, 962349563.3, 
    962349564.3, 962349565.3, 962349566.3, 962349567.3, 962349568.3, 
    962349569.3, 962349570.3, 962349571.3, 962349572.3, 962349572.8, 
    962349573.8, 962349574.8, 962349575.8, 962349576.8, 962349577.8, 
    962349578.8, 962349579.8, 962349580.8, 962349581.8, 962349582.8, 
    962349583.8, 962349584.8, 962349585.8, 962349586.8, 962349587.8, 
    962349588.8, 962349589.8, 962349590.8, 962349591.8, 962349592.8, 
    962349593.8, 962349594.8, 962349595.8, 962349596.8, 962349597.8, 
    962349598.8, 962349599.8, 962349600.8, 962349601.8, 962349602.8, 
    962349603.8, 962349604.8, 962349605.8, 962349606.8, 962349607.8, 
    962349608.8, 962349609.8, 962349610.8, 962349611.8, 962349612.8, 
    962349613.8, 962349614.3, 962349615.3, 962349616.3, 962349617.3, 
    962349618.3, 962349619.3, 962349620.3, 962349621.3, 962349622.3, 
    962349623.3, 962349623.8, 962349624.8, 962349625.8, 962349626.8, 
    962349627.8, 962349628.8, 962349629.8, 962349630.8, 962349631.8, 
    962349632.8, 962349633.8, 962349634.3, 962349635.3, 962349636.3, 
    962349637.3, 962349638.3, 962349639.3, 962349640.3, 962349641.3, 
    962349642.3, 962349642.8, 962349643.8, 962349644.4, 962349645.4, 
    962349646.4, 962349647.4, 962349648.4, 962349649.4, 962349650.4, 
    962349651.4, 962349652.4, 962349653.4, 962349654.4, 962349655.4, 
    962349656.4, 962349657.4, 962349658.4, 962349659.4, 962349660.4, 
    962349661.4, 962349662.4, 962349663.4, 962349664.4, 962349665.4, 
    962349666.4, 962349667.4, 962349668.4, 962349669.4, 962349670.4, 
    962349671.4, 962349672.4, 962349673.4, 962349674.4, 962349674.9, 
    962349675.9, 962349676.9, 962349677.9, 962349678.9, 962349679.9, 
    962349680.9, 962349681.9, 962349682.9, 962349683.9, 962349684.9, 
    962349685.9, 962349686.9, 962349687.9, 962349688.9, 962349689.9, 
    962349690.9, 962349691.9, 962349692.9, 962349693.9, 962349694.9, 
    962349695.9, 962349696.9, 962349697.9, 962349698.9, 962349699.9, 
    962349700.9, 962349701.9, 962349702.9, 962349703.9, 962349704.9, 
    962349705.9, 962349706.9, 962349707.9, 962349708.9, 962349709.9, 
    962349710.9, 962349711.9, 962349712.9, 962349713.9, 962349714.9, 
    962349715.4, 962349716.4, 962349717.4, 962349718.4, 962349719.4, 
    962349720.4, 962349721.4, 962349722.4, 962349723.4, 962349724.4, 
    962349725.4, 962349726.4, 962349727.4, 962349728.4, 962349729.4, 
    962349730.4, 962349731.4, 962349732.4, 962349733.4, 962349734.4, 
    962349735.5, 962349736.5, 962349737.5, 962349738.5, 962349739.5, 
    962349740.5, 962349741.5, 962349742.5, 962349743.5, 962349744.5, 
    962349745.5, 962349746.5, 962349747.5, 962349748.5, 962349749.5, 
    962349750.5, 962349751.5, 962349752.5, 962349753.5, 962349754.5, 
    962349755.5, 962349756.5, 962349757, 962349758, 962349759, 962349760, 
    962349761, 962349762, 962349763, 962349764, 962349765, 962349766, 
    962349767, 962349768, 962349769, 962349770, 962349771, 962349772, 
    962349773, 962349774, 962349775, 962349776, 962349777, 962349778, 
    962349779, 962349780, 962349781, 962349782, 962349783, 962349784, 
    962349785, 962349786, 962349787, 962349788, 962349789, 962349790, 
    962349791, 962349792, 962349793, 962349794, 962349795, 962349796, 
    962349797, 962349798, 962349798.5, 962349799.5, 962349800.5, 962349801.5, 
    962349802.5, 962349803.5, 962349804.5, 962349805.5, 962349806.5, 
    962349807.5, 962349808.5, 962349809.5, 962349810.5, 962349811.5, 
    962349812.5, 962349813.5, 962349814.5, 962349815.5, 962349816.5, 
    962349817.5, 962349818.5, 962349819.5, 962349820.5, 962349821.5, 
    962349822.5, 962349823.5, 962349824.5, 962349825.5, 962349826.5, 
    962349827.5, 962349828.5, 962349829.5, 962349830.5, 962349831.5, 
    962349832.5, 962349833.5, 962349834.5, 962349835.5, 962349836.5, 
    962349837.6, 962349838.6, 962349839.6, 962349840.6, 962349841.6, 
    962349842.6, 962349843.6, 962349844.6, 962349845.6, 962349846.6, 
    962349847.6, 962349848.6, 962349849.1, 962349850.1, 962349851.1, 
    962349852.1, 962349853.1, 962349854.1, 962349855.1, 962349856.1, 
    962349857.1, 962349858.1, 962349859.1, 962349860.1, 962349861.1, 
    962349862.1, 962349863.1, 962349864.1, 962349865.1, 962349866.1, 
    962349867.1, 962349868.1, 962349869.1, 962349870.1, 962349871.1, 
    962349872.1, 962349873.1, 962349874.1, 962349875.1, 962349876.1, 
    962349877.1, 962349878.1, 962349879.1, 962349880.1, 962349881.1, 
    962349882.1, 962349883.1, 962349884.1, 962349885.1, 962349886.1, 
    962349887.1, 962349888.1, 962349889.1, 962349890.1, 962349891.1, 
    962349892.1, 962349893.1, 962349894.1, 962349895.1, 962349896.1, 
    962349897.1, 962349898.1, 962349899.1, 962349899.6, 962349900.6, 
    962349901.6, 962349902.6, 962349903.6, 962349904.6, 962349905.6, 
    962349906.6, 962349907.6, 962349908.6, 962349909.6, 962349910.6, 
    962349911.6, 962349912.6, 962349913.6, 962349914.6, 962349915.6, 
    962349916.6, 962349917.6, 962349918.6, 962349919.6, 962349920.1, 
    962349921.1, 962349922.1, 962349923.1, 962349924.1, 962349925.1, 
    962349926.1, 962349927.1, 962349928.1, 962349929.1, 962349930.1, 
    962349931.1, 962349932.1, 962349933.1, 962349934.1, 962349935.1, 
    962349936.1, 962349937.1, 962349938.1, 962349939.1, 962349940.1, 
    962349941.1, 962349942.1, 962349943.1, 962349944.1, 962349945.1, 
    962349946.1, 962349947.1, 962349948.1, 962349949.1, 962349950.2, 
    962349951.2, 962349952.2, 962349953.2, 962349954.2, 962349955.2, 
    962349956.2, 962349957.2, 962349958.2, 962349959.2, 962349960.2, 
    962349961.2, 962349962.2, 962349963.2, 962349964.2, 962349965.2, 
    962349966.2, 962349967.2, 962349968.2, 962349969.2, 962349970.2, 
    962349971.2, 962349971.7, 962349972.7, 962349973.7, 962349974.7, 
    962349975.7, 962349976.7, 962349977.7, 962349978.7, 962349979.7, 
    962349980.7, 962349981.7, 962349982.7, 962349983.7, 962349984.7, 
    962349985.7, 962349986.7, 962349987.7, 962349988.7, 962349989.7, 
    962349990.7, 962349991.7, 962349992.7, 962349993.7, 962349994.7, 
    962349995.7, 962349996.7, 962349997.7, 962349998.7, 962349999.7, 
    962350000.7, 962350001.7, 962350002.7, 962350003.2, 962350004.2, 
    962350005.2, 962350006.2, 962350007.2, 962350008.2, 962350009.2, 
    962350010.2, 962350011.2, 962350011.7, 962350012.7, 962350013.7, 
    962350014.7, 962350015.7, 962350016.7, 962350017.7, 962350018.7, 
    962350019.7, 962350020.7, 962350021.7, 962350022.2, 962350023.2, 
    962350024.2, 962350025.2, 962350026.2, 962350027.2, 962350028.2, 
    962350029.2, 962350030.2, 962350031.2, 962350032.2, 962350032.7, 
    962350033.7, 962350034.7, 962350035.7, 962350036.7, 962350037.7, 
    962350038.7, 962350039.7, 962350040.7, 962350041.8, 962350042.8, 
    962350043.8, 962350044.8, 962350045.8, 962350046.8, 962350047.8, 
    962350048.8, 962350049.8, 962350050.8, 962350051.8, 962350052.8, 
    962350053.3, 962350054.3, 962350055.3, 962350056.3, 962350057.3, 
    962350058.3, 962350059.3, 962350060.3, 962350061.3, 962350062.3, 
    962350063.3, 962350063.8, 962350064.8, 962350065.8, 962350066.8, 
    962350067.8, 962350068.8, 962350069.8, 962350070.8, 962350071.8, 
    962350072.8, 962350073.8, 962350074.3, 962350075.3, 962350076.3, 
    962350077.3, 962350078.3, 962350079.3, 962350080.3, 962350081.3, 
    962350082.3, 962350083.3, 962350083.8, 962350084.8, 962350085.8, 
    962350086.8, 962350087.8, 962350088.8, 962350089.8, 962350090.8, 
    962350091.8, 962350092.8, 962350093.8, 962350094.8, 962350095.8, 
    962350096.8, 962350097.8, 962350098.8, 962350099.8, 962350100.8, 
    962350101.8, 962350102.8, 962350103.8, 962350104.3, 962350105.3, 
    962350106.3, 962350107.3, 962350108.3, 962350109.3, 962350110.3, 
    962350111.3, 962350112.3, 962350113.3, 962350114.3, 962350115.3, 
    962350116.3, 962350117.3, 962350118.3, 962350119.3, 962350120.3, 
    962350121.3, 962350122.3, 962350123.3, 962350124.3, 962350125.3, 
    962350126.3, 962350127.3, 962350128.3, 962350129.3, 962350130.3, 
    962350131.3, 962350132.3, 962350133.3, 962350134.3, 962350134.8, 
    962350135.8, 962350136.8, 962350137.8, 962350138.8, 962350139.8, 
    962350140.8, 962350141.8, 962350142.8, 962350143.8, 962350144.3, 
    962350145.3, 962350146.3, 962350147.3, 962350148.3, 962350149.3, 
    962350150.3, 962350151.3, 962350152.3, 962350153.3, 962350154.4, 
    962350155.4, 962350156.4, 962350157.4, 962350158.4, 962350159.4, 
    962350160.4, 962350161.4, 962350162.4, 962350163.4, 962350164.4, 
    962350164.9, 962350165.9, 962350166.9, 962350167.9, 962350168.9, 
    962350169.9, 962350170.9, 962350171.9, 962350172.9, 962350173.9, 
    962350174.9, 962350175.4, 962350176.4, 962350177.4, 962350178.4, 
    962350179.4, 962350180.4, 962350181.4, 962350182.4, 962350183.4, 
    962350184.4, 962350185.4, 962350185.9, 962350186.9, 962350187.9, 
    962350188.9, 962350189.9, 962350190.9, 962350191.9, 962350192.9, 
    962350193.9, 962350194.9, 962350195.9, 962350196.4, 962350197.4, 
    962350198.4, 962350199.4, 962350200.4, 962350201.4, 962350202.4, 
    962350203.4, 962350204.4, 962350205.4, 962350206.4, 962350206.9, 
    962350207.9, 962350208.9, 962350209.9, 962350210.9, 962350211.9, 
    962350212.9, 962350213.9, 962350214.9, 962350215.9, 962350216.9, 
    962350217.9, 962350218.9, 962350219.9, 962350220.9, 962350221.9, 
    962350222.9, 962350223.9, 962350224.9, 962350225.9, 962350226.9, 
    962350227.9, 962350228.9, 962350229.9, 962350230.9, 962350231.9, 
    962350232.9, 962350233.9, 962350234.9, 962350235.9, 962350236.9, 
    962350237.4, 962350238.4, 962350239.4, 962350240.4, 962350241.4, 
    962350242.4, 962350243.4, 962350244.4, 962350245.4, 962350246.5, 
    962350247.5, 962350248.5, 962350249.5, 962350250.5, 962350251.5, 
    962350252.5, 962350253.5, 962350254.5, 962350255.5, 962350256.5, 
    962350257, 962350258, 962350259, 962350260, 962350261, 962350262, 
    962350263, 962350264, 962350265, 962350266, 962350267, 962350268, 
    962350269, 962350270, 962350271, 962350272, 962350273, 962350274, 
    962350275, 962350276, 962350277, 962350277.5, 962350278.5, 962350279.5, 
    962350280.5, 962350281.5, 962350282.5, 962350283.5, 962350284.5, 
    962350285.5, 962350286.5, 962350287, 962350288, 962350289, 962350290, 
    962350291, 962350292, 962350293, 962350294, 962350295, 962350296, 
    962350297, 962350298, 962350298.5, 962350299.5, 962350300.5, 962350301.5, 
    962350302.5, 962350303.5, 962350304.5, 962350305.5, 962350306.5, 
    962350307.5, 962350308.5, 962350309.5, 962350310.5, 962350311.5, 
    962350312.5, 962350313.5, 962350314.5, 962350315.5, 962350316.5, 
    962350317.5, 962350318, 962350319, 962350320, 962350321, 962350322, 
    962350323, 962350324, 962350325, 962350326, 962350327, 962350328, 
    962350329, 962350329.5, 962350330.5, 962350331.5, 962350332.5, 
    962350333.5, 962350334.5, 962350335.5, 962350336.5, 962350337.5, 
    962350338.5, 962350339.5, 962350340.5, 962350341.5, 962350342.5, 
    962350343.5, 962350344.5, 962350345.5, 962350346.5, 962350347.5, 
    962350348.5, 962350349.1, 962350350.1, 962350351.1, 962350352.1, 
    962350353.1, 962350354.1, 962350355.1, 962350356.1, 962350357.1, 
    962350358.1, 962350358.6, 962350359.6, 962350360.6, 962350361.6, 
    962350362.6, 962350363.6, 962350364.6, 962350365.6, 962350366.6, 
    962350367.6, 962350368.6, 962350369.6, 962350370.6, 962350371.6, 
    962350372.6, 962350373.6, 962350374.6, 962350375.6, 962350376.6, 
    962350377.6, 962350378.6, 962350379.1, 962350380.1, 962350381.1, 
    962350382.1, 962350383.1, 962350384.1, 962350385.1, 962350386.1, 
    962350387.1, 962350388.1, 962350389.1, 962350390.1, 962350391.1, 
    962350392.1, 962350393.1, 962350394.1, 962350395.1, 962350396.1, 
    962350397.1, 962350398.1, 962350399.1, 962350400.1, 962350401.1, 
    962350402.1, 962350403.1, 962350404.1, 962350405.1, 962350406.1, 
    962350407.1, 962350408.1, 962350409.1, 962350410.1, 962350411.1, 
    962350411.6, 962350412.6, 962350413.6, 962350414.6, 962350415.6 ;
}
